module main(
a,
b,
out
);

	input a;
	input b;
	output out;

	and(out, a, b);



endmodule
